// Start Positions maps given STARTpos to set of pixels for display
module startPositions (STARTpos, PixSTART);
	input logic [3:0] STARTpos;
	output logic [15:0][15:0] PixSTART;
	
	always_comb begin
		case (STARTpos)
			0: PixSTART = '0;
			
			1: begin
				PixSTART[00] = 16'b0000000000000000;
				PixSTART[01] = 16'b0000000000000000;
				PixSTART[02] = 16'b0000000000000000;
				PixSTART[03] = 16'b0000001111000000;
				PixSTART[04] = 16'b0000010000100000;
				PixSTART[05] = 16'b0000000000100000;
				PixSTART[06] = 16'b0000000000100000;
				PixSTART[07] = 16'b0000000000100000;
				PixSTART[08] = 16'b0000000111000000;
				PixSTART[09] = 16'b0000000000100000;
				PixSTART[10] = 16'b0000000000100000;
				PixSTART[11] = 16'b0000010000100000;
				PixSTART[12] = 16'b0000001111000000;
				PixSTART[13] = 16'b0000000000000000;
				PixSTART[14] = 16'b0000000000000000;
				PixSTART[15] = 16'b0000000000000000;
			end
			
			2: begin
				PixSTART[00] = 16'b0000000000000000;
				PixSTART[01] = 16'b0000000000000000;
				PixSTART[02] = 16'b0000000000000000;
				PixSTART[03] = 16'b0000001111000000;
				PixSTART[04] = 16'b0000010000100000;
				PixSTART[05] = 16'b0000000000100000;
				PixSTART[06] = 16'b0000000000100000;
				PixSTART[07] = 16'b0000000001000000;
				PixSTART[08] = 16'b0000000010000000;
				PixSTART[09] = 16'b0000000100000000;
				PixSTART[10] = 16'b0000001000000000;
				PixSTART[11] = 16'b0000010000000000;
				PixSTART[12] = 16'b0000011111100000;
				PixSTART[13] = 16'b0000000000000000;
				PixSTART[14] = 16'b0000000000000000;
				PixSTART[15] = 16'b0000000000000000;
			end
			
			3: begin
				PixSTART[00] = 16'b0000000000000000;
				PixSTART[01] = 16'b0000000000000000;
				PixSTART[02] = 16'b0000000000000000;
				PixSTART[03] = 16'b0000001110000000;
				PixSTART[04] = 16'b0000010010000000;
				PixSTART[05] = 16'b0000000010000000;
				PixSTART[06] = 16'b0000000010000000;
				PixSTART[07] = 16'b0000000010000000;
				PixSTART[08] = 16'b0000000010000000;
				PixSTART[09] = 16'b0000000010000000;
				PixSTART[10] = 16'b0000000010000000;
				PixSTART[11] = 16'b0000000010000000;
				PixSTART[12] = 16'b0000001111000000;
				PixSTART[13] = 16'b0000000000000000;
				PixSTART[14] = 16'b0000000000000000;
				PixSTART[15] = 16'b0000000000000000;
			end
			
			default: begin
				PixSTART[00] = 16'b0000000000000000;
				PixSTART[01] = 16'b0000000000000000;
				PixSTART[02] = 16'b0000000000000000;
				PixSTART[03] = 16'b0111100011110011;
				PixSTART[04] = 16'b1000010100001011;
				PixSTART[05] = 16'b1000000100001011;
				PixSTART[06] = 16'b1000000100001011;
				PixSTART[07] = 16'b1000000100001011;
				PixSTART[08] = 16'b1000000100001011;
				PixSTART[09] = 16'b1001100100001011;
				PixSTART[10] = 16'b1000100100001000;
				PixSTART[11] = 16'b1000100100001011;
				PixSTART[12] = 16'b0111000011110011;
				PixSTART[13] = 16'b0000000000000000;
				PixSTART[14] = 16'b0000000000000000;
				PixSTART[15] = 16'b0000000000000000;
			end
		endcase
	end
endmodule