module endExplode (position, PixEND);
	input logic [3:0] position;
	output logic [15:0][15:0] PixEND;
	
	
	always_comb begin
		case (position)
			0: PixEND = '0;
			
			1: begin // Explode Position 0
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0000000000000000;
				PixEND[06] = 16'b0000000000000000;
				PixEND[07] = 16'b0000001100000000;
				PixEND[08] = 16'b0000001100000000;
				PixEND[09] = 16'b0000000000000000;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			2: begin // Explode Position 1
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0000100001000000;
				PixEND[06] = 16'b0000010010000000;
				PixEND[07] = 16'b0000001100000000;
				PixEND[08] = 16'b0000001100000000;
				PixEND[09] = 16'b0000010010000000;
				PixEND[10] = 16'b0000100001000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			3: begin // Explode Position 2
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0010001100010000;
				PixEND[04] = 16'b0001010010100000;
				PixEND[05] = 16'b0000100001000000;
				PixEND[06] = 16'b0000010010000000;
				PixEND[07] = 16'b0000001100000000;
				PixEND[08] = 16'b0000001100000000;
				PixEND[09] = 16'b0000010010000000;
				PixEND[10] = 16'b0000100001000000;
				PixEND[11] = 16'b0001010010100000;
				PixEND[12] = 16'b0010001100010000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			4: begin // Explode Position 3
				PixEND[00] = 16'b0001000010000000;
				PixEND[01] = 16'b0010000100000000;
				PixEND[02] = 16'b0100001000000000;
				PixEND[03] = 16'b0010001100010000;
				PixEND[04] = 16'b0001010010100000;
				PixEND[05] = 16'b0000100001010000;
				PixEND[06] = 16'b0000010010001000;
				PixEND[07] = 16'b0000001100000100;
				PixEND[08] = 16'b0000001100000000;
				PixEND[09] = 16'b0000010010000000;
				PixEND[10] = 16'b0000100001000000;
				PixEND[11] = 16'b0001010010100000;
				PixEND[12] = 16'b0010001100010000;
				PixEND[13] = 16'b0010000010000000;
				PixEND[14] = 16'b0001000001000000;
				PixEND[15] = 16'b0010000000000000;
			end
			
			5: begin // ALL RED
				PixEND = '1;
			end
			
			6: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			7: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			8: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			9: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			10: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			11: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			12: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			13: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			14: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			15: begin // END
				PixEND[00] = 16'b0000000000000000;
				PixEND[01] = 16'b0000000000000000;
				PixEND[02] = 16'b0000000000000000;
				PixEND[03] = 16'b0000000000000000;
				PixEND[04] = 16'b0000000000000000;
				PixEND[05] = 16'b0111010001011100;
				PixEND[06] = 16'b0100011001010010;
				PixEND[07] = 16'b0111010101010010;
				PixEND[08] = 16'b0100010011010010;
				PixEND[09] = 16'b0111010001011100;
				PixEND[10] = 16'b0000000000000000;
				PixEND[11] = 16'b0000000000000000;
				PixEND[12] = 16'b0000000000000000;
				PixEND[13] = 16'b0000000000000000;
				PixEND[14] = 16'b0000000000000000;
				PixEND[15] = 16'b0000000000000000;
			end
			
			default: PixEND = '0;
		endcase
	end
endmodule

//module endExplode_testbench();
//	logic [3:0]	position;
//	logic [15:0][15:0] PixEND;
//	
//	endExplode dut (.position, .PixEND);
//	
//	integer i;
//	initial begin
//		for (i=0; i<8; i++) begin
//			position = i; #10;
//		end
//	end
//endmodule