module collisionCheck (in, out);
	input logic [15:0][15:0] in;
	output logic out;
	
	assign out = in[00][00]|in[00][01]|in[00][02]|in[00][03]|in[00][04]|in[00][05]|in[00][06]|in[00][07]|in[00][08]|in[00][09]|in[00][10]|in[00][11]|in[00][12]|in[00][13]|in[00][14]|in[00][15]
					|in[01][00]|in[01][01]|in[01][02]|in[01][03]|in[01][04]|in[01][05]|in[01][06]|in[01][07]|in[01][08]|in[01][09]|in[01][10]|in[01][11]|in[01][12]|in[01][13]|in[01][14]|in[01][15]
					|in[02][00]|in[02][01]|in[02][02]|in[02][03]|in[02][04]|in[02][05]|in[02][06]|in[02][07]|in[02][08]|in[02][09]|in[02][10]|in[02][11]|in[02][12]|in[02][13]|in[02][14]|in[02][15]
					|in[03][00]|in[03][01]|in[03][02]|in[03][03]|in[03][04]|in[03][05]|in[03][06]|in[03][07]|in[03][08]|in[03][09]|in[03][10]|in[03][11]|in[03][12]|in[03][13]|in[03][14]|in[03][15]
					|in[04][00]|in[04][01]|in[04][02]|in[04][03]|in[04][04]|in[04][05]|in[04][06]|in[04][07]|in[04][08]|in[04][09]|in[04][10]|in[04][11]|in[04][12]|in[04][13]|in[04][14]|in[04][15]
					|in[05][00]|in[05][01]|in[05][02]|in[05][03]|in[05][04]|in[05][05]|in[05][06]|in[05][07]|in[05][08]|in[05][09]|in[05][10]|in[05][11]|in[05][12]|in[05][13]|in[05][14]|in[05][15]
					|in[06][00]|in[06][01]|in[06][02]|in[06][03]|in[06][04]|in[06][05]|in[06][06]|in[06][07]|in[06][08]|in[06][09]|in[06][10]|in[06][11]|in[06][12]|in[06][13]|in[06][14]|in[06][15]
					|in[07][00]|in[07][01]|in[07][02]|in[07][03]|in[07][04]|in[07][05]|in[07][06]|in[07][07]|in[07][08]|in[07][09]|in[07][10]|in[07][11]|in[07][12]|in[07][13]|in[07][14]|in[07][15]
					|in[08][00]|in[08][01]|in[08][02]|in[08][03]|in[08][04]|in[08][05]|in[08][06]|in[08][07]|in[08][08]|in[08][09]|in[08][10]|in[08][11]|in[08][12]|in[08][13]|in[08][14]|in[08][15]
					|in[09][00]|in[09][01]|in[09][02]|in[09][03]|in[09][04]|in[09][05]|in[09][06]|in[09][07]|in[09][08]|in[09][09]|in[09][10]|in[09][11]|in[09][12]|in[09][13]|in[09][14]|in[09][15]
					|in[10][00]|in[10][01]|in[10][02]|in[10][03]|in[10][04]|in[10][05]|in[10][06]|in[10][07]|in[10][08]|in[10][09]|in[10][10]|in[10][11]|in[10][12]|in[10][13]|in[10][14]|in[10][15]
					|in[11][00]|in[11][01]|in[11][02]|in[11][03]|in[11][04]|in[11][05]|in[11][06]|in[11][07]|in[11][08]|in[11][09]|in[11][10]|in[11][11]|in[11][12]|in[11][13]|in[11][14]|in[11][15]
					|in[12][00]|in[12][01]|in[12][02]|in[12][03]|in[12][04]|in[12][05]|in[12][06]|in[12][07]|in[12][08]|in[12][09]|in[12][10]|in[12][11]|in[12][12]|in[12][13]|in[12][14]|in[12][15]
					|in[13][00]|in[13][01]|in[13][02]|in[13][03]|in[13][04]|in[13][05]|in[13][06]|in[13][07]|in[13][08]|in[13][09]|in[13][10]|in[13][11]|in[13][12]|in[13][13]|in[13][14]|in[13][15]
					|in[14][00]|in[14][01]|in[14][02]|in[14][03]|in[14][04]|in[14][05]|in[14][06]|in[14][07]|in[14][08]|in[14][09]|in[14][10]|in[14][11]|in[14][12]|in[14][13]|in[14][14]|in[14][15]
					|in[15][00]|in[15][01]|in[15][02]|in[15][03]|in[15][04]|in[15][05]|in[15][06]|in[15][07]|in[15][08]|in[15][09]|in[15][10]|in[15][11]|in[15][12]|in[15][13]|in[15][14]|in[15][15];
endmodule

//module collisionCheck_testbench();
//	logic out;
//	logic [15:0][15:0] in;
//	
//	collisionCheck dut (.in, .out);
//	
//	initial begin
//		in <= '0; #10;
//		in[5][14] <= 1; #10;
//		in <= '0; #10;
//		in[0][0] <= 1; #10;
//	end
//endmodule